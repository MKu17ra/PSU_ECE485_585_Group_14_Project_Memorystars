
`timescale 1ns/1ns

module tb();
	initial begin
		$display("ece585 - Julia Filipchuk");
	end
endmodule : tb

